----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03.02.2022 17:51:12
-- Design Name: 
-- Module Name: ModuloDEC - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ModuloDEC is
    Port ( S : in STD_LOGIC_VECTOR (3 downto 0);
           O : out STD_LOGIC_VECTOR (6 downto 0));
end ModuloDEC;

architecture Behavioral of ModuloDEC is

begin

with S select 
    O <= "0000001" when "0000",
         "1001111" when "0001",
         "0010010" when "0010",
         "0000110" when "0011",
         "1001100" when "0100",
         "0100100" when "0101",
         "1100000" when "0110",
         "0001110" when "0111",
         "0000000" when "1000",
         "0000100" when "1001",
         "1111110" when "1010",
         "0110000" when "1011",
         "1101101" when "1100",
         "1111001" when "1101",
         "0110011" when "1110",
         "1011011" when others;

end Behavioral;
